--------------------------------------------------------------------------------
-- Project :
-- File    :
-- Autor   :
-- Date    :
--
--------------------------------------------------------------------------------
-- Description :
--
--------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Reg_file IS
  PORT (
    clock,write_e, reset      : IN  std_logic;
    rd1a,rd2a,rwa,manual_address : IN std_logic_vector(4 DOWNTO 0);
    rw : IN std_logic_vector (31 DOWNTO 0);

    rd1,rd2, manual_value        : OUT std_logic_vector(31 DOWNTO 0)
    );
END Reg_file;

--------------------------------------------------------------------------------
--Complete your VHDL description below
--------------------------------------------------------------------------------

ARCHITECTURE TypeArchitecture OF Reg_file IS
TYPE register_file is array(0 to 31) of std_logic_vector(31 DOWNTO 0);
SIGNAL registers : register_file := 
   ("00000000000000000000000000000000","00000000000000000000000000001000","00000000000000000000000000000010","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000");
BEGIN
process (clock, write_e, reset, registers, rd1a, rd2a, rwa, rw, manual_address)
BEGIN
manual_value <= registers(to_integer(unsigned(manual_address)));
IF (1 = 1) THEN
	rd1 <= registers(to_integer(unsigned(rd1a)));
	rd2 <= registers(to_integer(unsigned(rd2a)));
	IF (write_e = '1' AND to_integer(unsigned(rwa)) /= 0) THEN --Can't write on register X0
		registers(to_integer(unsigned(rwa))) <= rw;
	END IF;
END IF;
IF (reset = '1') THEN --Wipes all registers
	registers <= 
   ("00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000");
END IF;
END PROCESS;
END TypeArchitecture;
