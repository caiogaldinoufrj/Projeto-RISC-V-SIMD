--------------------------------------------------------------------------------
-- Project :
-- File    :
-- Autor   :
-- Date    :
--
--------------------------------------------------------------------------------
-- Description :
--
--------------------------------------------------------------------------------

library IEEE;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

 entity Somador is

  port(A, B_u : in std_logic_vector (31 downto 0);
  S : out std_logic_vector (31 downto 0));

 end Somador;

 architecture TypeArchitecture of Somador is
 signal C     : std_logic_vector (31 downto 0);
 signal control  : std_logic_vector (2 downto 0);
 signal mode : std_logic;
 begin
 
    control(0) <= '1';
    control(1) <= '1';
    control(2) <= '1';
    mode <= '0';
    
Carrys:process(C, control, mode, A, B_u)
begin
    C(0) <= mode;
    C(1) <= (A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode));
    C(2) <= (A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))));
    C(3) <= (A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))));
    C(4) <= (((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)));
    C(5) <= (A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))));
    C(6) <= (A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))));
    C(7) <= (A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))));
    C(8) <= (((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)));
    C(9) <= (A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))));
    C(10) <= (A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))));
    C(11) <= (A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))));
    C(12) <= (((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)));
    C(13) <= (A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))));
    C(14) <= (A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))));
    C(15) <= (A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))));
    C(16) <= (((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)));
    C(17) <= (A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))));
    C(18) <= (A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))));
    C(19) <= (A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))));
    C(20) <= (((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)));
    C(21) <= (A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))));
    C(22) <= (A(21) and B_u(21)) or ((A(21) or B_u(21)) and ((A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))))));
    C(23) <= (A(22) and B_u(22)) or ((A(22) or B_u(22)) and ((A(21) and B_u(21)) or ((A(21) or B_u(21)) and ((A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))))))));
    C(24) <= (((A(23) and B_u(23)) or ((A(23) or B_u(23)) and ((A(22) and B_u(22)) or ((A(22) or B_u(22)) and ((A(21) and B_u(21)) or ((A(21) or B_u(21)) and ((A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)));
    C(25) <= (A(24) and B_u(24)) or ((A(24) or B_u(24)) and ((((A(23) and B_u(23)) or ((A(23) or B_u(23)) and ((A(22) and B_u(22)) or ((A(22) or B_u(22)) and ((A(21) and B_u(21)) or ((A(21) or B_u(21)) and ((A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))));
    C(26) <= (A(25) and B_u(25)) or ((A(25) or B_u(25)) and ((A(24) and B_u(24)) or ((A(24) or B_u(24)) and ((((A(23) and B_u(23)) or ((A(23) or B_u(23)) and ((A(22) and B_u(22)) or ((A(22) or B_u(22)) and ((A(21) and B_u(21)) or ((A(21) or B_u(21)) and ((A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))));
    C(27) <= (A(26) and B_u(26)) or ((A(26) or B_u(26)) and ((A(25) and B_u(25)) or ((A(25) or B_u(25)) and ((A(24) and B_u(24)) or ((A(24) or B_u(24)) and ((((A(23) and B_u(23)) or ((A(23) or B_u(23)) and ((A(22) and B_u(22)) or ((A(22) or B_u(22)) and ((A(21) and B_u(21)) or ((A(21) or B_u(21)) and ((A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))));
    C(28) <= (((A(27) and B_u(27)) or ((A(27) or B_u(27)) and ((A(26) and B_u(26)) or ((A(26) or B_u(26)) and ((A(25) and B_u(25)) or ((A(25) or B_u(25)) and ((A(24) and B_u(24)) or ((A(24) or B_u(24)) and ((((A(23) and B_u(23)) or ((A(23) or B_u(23)) and ((A(22) and B_u(22)) or ((A(22) or B_u(22)) and ((A(21) and B_u(21)) or ((A(21) or B_u(21)) and ((A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)));
    C(29) <= (A(28) and B_u(28)) or ((A(28) or B_u(28)) and ((((A(27) and B_u(27)) or ((A(27) or B_u(27)) and ((A(26) and B_u(26)) or ((A(26) or B_u(26)) and ((A(25) and B_u(25)) or ((A(25) or B_u(25)) and ((A(24) and B_u(24)) or ((A(24) or B_u(24)) and ((((A(23) and B_u(23)) or ((A(23) or B_u(23)) and ((A(22) and B_u(22)) or ((A(22) or B_u(22)) and ((A(21) and B_u(21)) or ((A(21) or B_u(21)) and ((A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))));
    C(30) <= (A(29) and B_u(29)) or ((A(29) or B_u(29)) and ((A(28) and B_u(28)) or ((A(28) or B_u(28)) and ((((A(27) and B_u(27)) or ((A(27) or B_u(27)) and ((A(26) and B_u(26)) or ((A(26) or B_u(26)) and ((A(25) and B_u(25)) or ((A(25) or B_u(25)) and ((A(24) and B_u(24)) or ((A(24) or B_u(24)) and ((((A(23) and B_u(23)) or ((A(23) or B_u(23)) and ((A(22) and B_u(22)) or ((A(22) or B_u(22)) and ((A(21) and B_u(21)) or ((A(21) or B_u(21)) and ((A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))));
    C(31) <= (A(30) and B_u(30)) or ((A(30) or B_u(30)) and ((A(29) and B_u(29)) or ((A(29) or B_u(29)) and ((A(28) and B_u(28)) or ((A(28) or B_u(28)) and ((((A(27) and B_u(27)) or ((A(27) or B_u(27)) and ((A(26) and B_u(26)) or ((A(26) or B_u(26)) and ((A(25) and B_u(25)) or ((A(25) or B_u(25)) and ((A(24) and B_u(24)) or ((A(24) or B_u(24)) and ((((A(23) and B_u(23)) or ((A(23) or B_u(23)) and ((A(22) and B_u(22)) or ((A(22) or B_u(22)) and ((A(21) and B_u(21)) or ((A(21) or B_u(21)) and ((A(20) and B_u(20)) or ((A(20) or B_u(20)) and ((((A(19) and B_u(19)) or ((A(19) or B_u(19)) and ((A(18) and B_u(18)) or ((A(18) or B_u(18)) and ((A(17) and B_u(17)) or ((A(17) or B_u(17)) and ((A(16) and B_u(16)) or ((A(16) or B_u(16)) and ((((A(15) and B_u(15)) or ((A(15) or B_u(15)) and ((A(14) and B_u(14)) or ((A(14) or B_u(14)) and ((A(13) and B_u(13)) or ((A(13) or B_u(13)) and ((A(12) and B_u(12)) or ((A(12) or B_u(12)) and ((((A(11) and B_u(11)) or ((A(11) or B_u(11)) and ((A(10) and B_u(10)) or ((A(10) or B_u(10)) and ((A(9) and B_u(9)) or ((A(9) or B_u(9)) and ((A(8) and B_u(8)) or ((A(8) or B_u(8)) and ((((A(7) and B_u(7)) or ((A(7) or B_u(7)) and ((A(6) and B_u(6)) or ((A(6) or B_u(6)) and ((A(5) and B_u(5)) or ((A(5) or B_u(5)) and ((A(4) and B_u(4)) or ((A(4) or B_u(4)) and ((((A(3) and B_u(3)) or ((A(3) or B_u(3)) and ((A(2) and B_u(2)) or ((A(2) or B_u(2)) and ((A(1) and B_u(1)) or ((A(1) or B_u(1)) and ((A(0) and B_u(0)) or ((A(0) or B_u(0)) and (mode))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(2)) or (mode and (not control(2)))))))))))) and control(0)) or (mode and (not control(0)))))))))))) and control(1)) or (mode and (not control(1)))))))))))) and control(0)) or (mode and (not control(0)))))))));

end process Carrys;
process(A,B_u,C)
    begin
    for n in 0 to 31 loop
      S(n) <= (A(n)xor B_u(n)) xor C(n);
    end loop;
    end process;
end TypeArchitecture;
